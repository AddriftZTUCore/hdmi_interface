`ifndef __TOP_DEFINE_VH
`define __TOP_DEFINE_VH 1

`define rst_block posedge clk or negedge rst_n
`define rst       !rst_n
`define RST_POSITIVE 0

`define FPGA_K7

`endif
